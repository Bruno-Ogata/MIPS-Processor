module Hard_Disk (
    input Clock,
	 //input [3:0] indice,            // Índice do programa (4 bits para até 10 programas)
    input [11:0] addr,              // Endereço dentro do programa
    output reg [31:0] instrucao    // Instrução lida
);
    reg [31:0] memoria_hd [0:2047]; // Memória total do HD (10 programas de 102 instruções)

    initial begin
        // Carregue os programas aqui
        // Exemplo: memória_hd[0] a memória_hd[99] -> Programa 0
        // memória_hd[100] a memória_hd[199] -> Programa 1, e assim por diante
		  
		  // Teste - Media 
		  memoria_hd[0] = 32'b00011100000000000000000000000001; // jump 1  
		  memoria_hd[1] = 32'b00000100000111010000000000101000; // addi $fp $zero 40
		  memoria_hd[2] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[3] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[4] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[5] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[6] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[7] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[8] = 32'b00101100000000101111111111111111; // input $t2
		  memoria_hd[9] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[10] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[11] = 32'b00001111101000110000000000000001; // lw $fp $t3 1
		  memoria_hd[12] = 32'b00101100000001001111111111111111; // input $t4
		  memoria_hd[13] = 32'b00000100100000110000000000000000; // addi $t3 $t4 0
		  memoria_hd[14] = 32'b00010011101000110000000000000001; // sw $fp $t3 1
		  memoria_hd[15] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[16] = 32'b00101100000001101111111111111111; // input $t6
		  memoria_hd[17] = 32'b00000100110001010000000000000000; // addi $t5 $t6 0
		  memoria_hd[18] = 32'b00010011101001010000000000000010; // sw $fp $t5 2
		  memoria_hd[19] = 32'b00001111101001110000000000000011; // lw $fp $t7 3
		  memoria_hd[20] = 32'b00001111101010000000000000000000; // lw $fp $t8 0
		  memoria_hd[21] = 32'b00001111101010010000000000000001; // lw $fp $t9 1
		  memoria_hd[22] = 32'b00000001000010010101000000000000; // add $t10 $t8 $t9
		  memoria_hd[23] = 32'b00001111101010110000000000000010; // lw $fp $t11 2
		  memoria_hd[24] = 32'b00000001010010110110000000000000; // add $t12 $t10 $t11
		  memoria_hd[25] = 32'b00000100000110110000000000000011; // addi $aux $zero 3
		  memoria_hd[26] = 32'b00000001100110110110100000000011; // div $t13 $t12 $aux
		  memoria_hd[27] = 32'b00000101101001110000000000000000; // addi $t7 $t13 0
		  memoria_hd[28] = 32'b00010011101001110000000000000011; // sw $fp $t7 3
		  memoria_hd[29] = 32'b00001111101011100000000000000011; // lw $fp $t14 3
		  memoria_hd[30] = 32'b00101001110111111111111111111111; // output $t14
		  memoria_hd[31] = 32'b11111000000000000000000000000000; // halt
		  
		  // Programa 1 - GCD
		  memoria_hd[200] = 32'b00011100000000000000000001001101; // jump 77
		  memoria_hd[201] = 32'b00010011101111110000000000000001; // sw $fp $ra 1
		  memoria_hd[202] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[203] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[204] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[205] = 32'b00001111101000010000000000000010; // lw $fp $t1 2
		  memoria_hd[206] = 32'b00001111101000100000000000000011; // lw $fp $t2 3
		  memoria_hd[207] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[208] = 32'b00001111101001000000000000000100; // lw $fp $t4 4
		  memoria_hd[209] = 32'b00000100100001000000000000000000; // addi $t4 $t4 0
		  memoria_hd[210] = 32'b00010011101001000000000000000100; // sw $fp $t4 4
		  memoria_hd[211] = 32'b00000000001000100010100000100101; // sge $t5 $t1 $t2
		  memoria_hd[212] = 32'b00010100000001010000000000011011; // beq $t5 $zero 27
		  memoria_hd[213] = 32'b00001111101001100000000000000010; // lw $fp $t6 2
		  memoria_hd[214] = 32'b00001111101001110000000000000010; // lw $fp $t7 2
		  memoria_hd[215] = 32'b00001111101010000000000000000011; // lw $fp $t8 3
		  memoria_hd[216] = 32'b00000000111010000100100000000001; // sub $t9 $t7 $t8
		  memoria_hd[217] = 32'b00000101001001100000000000000000; // addi $t6 $t9 0
		  memoria_hd[218] = 32'b00010011101001100000000000000010; // sw $fp $t6 2
		  memoria_hd[219] = 32'b00001111101010100000000000000100; // lw $fp $t10 4
		  memoria_hd[220] = 32'b00001111101010110000000000000100; // lw $fp $t11 4
		  memoria_hd[221] = 32'b00000100000110110000000000000001; // addi $aux $zero 1
		  memoria_hd[222] = 32'b00000001011110110110000000000000; // add $t12 $t11 $aux
		  memoria_hd[223] = 32'b00000101100010100000000000000000; // addi $t10 $t12 0
		  memoria_hd[224] = 32'b00010011101010100000000000000100; // sw $fp $t10 4
		  memoria_hd[225] = 32'b00000101100000010000000000000000; // addi $t1 $t12 0
		  memoria_hd[226] = 32'b00011100000000000000000000001011; // jump 11
		  memoria_hd[227] = 32'b00001111101011010000000000000100; // lw $fp $t13 4
		  memoria_hd[228] = 32'b00000101101111000000000000000000; // addi $gp $t13 0
		  memoria_hd[229] = 32'b00001111101111110000000000000001; // lw $fp $ra 1
		  memoria_hd[230] = 32'b00100111111000000000000000000000; // jr $ra $zero $zero
		  memoria_hd[231] = 32'b00010011101111110000000000000001; // sw $fp $ra 1
		  memoria_hd[232] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[233] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[234] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[235] = 32'b00001111101000010000000000000010; // lw $fp $t1 2
		  memoria_hd[236] = 32'b00001111101000100000000000000011; // lw $fp $t2 3
		  memoria_hd[237] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[238] = 32'b00000100000110110000000000000000; // addi $aux $zero 0
		  memoria_hd[239] = 32'b00000000010110110010000000000001; // sub $t4 $t2 $aux
		  memoria_hd[240] = 32'b00011000000001000000000000101100; // bne $t4 $zero 44
		  memoria_hd[241] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[242] = 32'b00000100101111000000000000000000; // addi $gp $t5 0
		  memoria_hd[243] = 32'b00011100000000000000000001001011; // jump 75
		  memoria_hd[244] = 32'b00001111101001100000000000000100; // lw $fp $t6 4
		  memoria_hd[245] = 32'b00001111101001110000000000000010; // lw $fp $t7 2
		  memoria_hd[246] = 32'b00001111101010000000000000000011; // lw $fp $t8 3
		  memoria_hd[247] = 32'b00010011110111010000000000000000; // sw $sp $fp 0
		  memoria_hd[248] = 32'b00000111110111010000000000000000; // addi $fp $sp 0
		  memoria_hd[249] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[250] = 32'b00010011101010000000000000000011; // sw $fp $t8 3
		  memoria_hd[251] = 32'b00010011101001110000000000000010; // sw $fp $t7 2
		  memoria_hd[252] = 32'b00110000000000000000000000000001; // jal 1
		  memoria_hd[253] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[254] = 32'b00001111101111010000000000000000; // lw $fp $fp 0
		  memoria_hd[255] = 32'b00000111100010010000000000000000; // addi $t9 $gp 0
		  memoria_hd[256] = 32'b00000101001001100000000000000000; // addi $t6 $t9 0
		  memoria_hd[257] = 32'b00010011101001100000000000000100; // sw $fp $t6 4
		  memoria_hd[258] = 32'b00001111101010100000000000000011; // lw $fp $t10 3
		  memoria_hd[259] = 32'b00001111101010110000000000000010; // lw $fp $t11 2
		  memoria_hd[260] = 32'b00001111101011000000000000000011; // lw $fp $t12 3
		  memoria_hd[261] = 32'b00001111101011010000000000000100; // lw $fp $t13 4
		  memoria_hd[262] = 32'b00000001100011010111000000000010; // mult $t14 $t12 $t13
		  memoria_hd[263] = 32'b00000001011011100111100000000001; // sub $t15 $t11 $t14
		  memoria_hd[264] = 32'b00010011110111010000000000000000; // sw $sp $fp 0
		  memoria_hd[265] = 32'b00000111110111010000000000000000; // addi $fp $sp 0
		  memoria_hd[266] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[267] = 32'b00010011101011110000000000000011; // sw $fp $t15 3
		  memoria_hd[268] = 32'b00010011101010100000000000000010; // sw $fp $t10 2
		  memoria_hd[269] = 32'b00110000000000000000000000011111; // jal 31
		  memoria_hd[270] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[271] = 32'b00001111101111010000000000000000; // lw $fp $fp 0
		  memoria_hd[272] = 32'b00000111100100000000000000000000; // addi $t16 $gp 0
		  memoria_hd[273] = 32'b00000110000111000000000000000000; // addi $gp $t16 0
		  memoria_hd[274] = 32'b00011100000000000000000001001011; // jump 75
		  memoria_hd[275] = 32'b00001111101111110000000000000001; // lw $fp $ra 1
		  memoria_hd[276] = 32'b00100111111000000000000000000000; // jr $ra $zero $zero
		  memoria_hd[277] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[278] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[279] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[280] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[281] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[282] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[283] = 32'b00101100000000101111111111111111; // input $t2
		  memoria_hd[284] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[285] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[286] = 32'b00001111101000110000000000000001; // lw $fp $t3 1
		  memoria_hd[287] = 32'b00101100000001001111111111111111; // input $t4
		  memoria_hd[288] = 32'b00000100100000110000000000000000; // addi $t3 $t4 0
		  memoria_hd[289] = 32'b00010011101000110000000000000001; // sw $fp $t3 1
		  memoria_hd[290] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[291] = 32'b00001111101001100000000000000000; // lw $fp $t6 0
		  memoria_hd[292] = 32'b00001111101001110000000000000001; // lw $fp $t7 1
		  memoria_hd[293] = 32'b00010011110111010000000000000000; // sw $sp $fp 0
		  memoria_hd[294] = 32'b00000111110111010000000000000000; // addi $fp $sp 0
		  memoria_hd[295] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[296] = 32'b00010011101001110000000000000011; // sw $fp $t7 3
		  memoria_hd[297] = 32'b00010011101001100000000000000010; // sw $fp $t6 2
		  memoria_hd[298] = 32'b00110000000000000000000000011111; // jal 31
		  memoria_hd[299] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[300] = 32'b00001111101111010000000000000000; // lw $fp $fp 0
		  memoria_hd[301] = 32'b00000111100010000000000000000000; // addi $t8 $gp 0
		  memoria_hd[302] = 32'b00000101000001010000000000000000; // addi $t5 $t8 0
		  memoria_hd[303] = 32'b00010011101001010000000000000010; // sw $fp $t5 2
		  memoria_hd[304] = 32'b00001111101010010000000000000010; // lw $fp $t9 2
		  memoria_hd[305] = 32'b00101001001111111111111111111111; // output $t9
		  memoria_hd[306] = 32'b11111000000000000000000000000000; // halt 
		  
		  // Programa 2 - Fibonacci 
		  memoria_hd[350] = 32'b00011100000000000000000000111000; // jump 56
		  memoria_hd[351] = 32'b00010011101111110000000000000001; // sw $fp $ra 1
		  memoria_hd[352] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[353] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[354] = 32'b00001111101000010000000000000010; // lw $fp $t1 2
		  memoria_hd[355] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[356] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[357] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[358] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[359] = 32'b00001111101000110000000000000011; // lw $fp $t3 3
		  memoria_hd[360] = 32'b00000100011000110000000000000000; // addi $t3 $t3 0
		  memoria_hd[361] = 32'b00010011101000110000000000000011; // sw $fp $t3 3
		  memoria_hd[362] = 32'b00001111101001000000000000000100; // lw $fp $t4 4
		  memoria_hd[363] = 32'b00000100100001000000000000000001; // addi $t4 $t4 1
		  memoria_hd[364] = 32'b00010011101001000000000000000100; // sw $fp $t4 4
		  memoria_hd[365] = 32'b00001111101001010000000000000110; // lw $fp $t5 6
		  memoria_hd[366] = 32'b00000100101001010000000000000010; // addi $t5 $t5 2
		  memoria_hd[367] = 32'b00010011101001010000000000000110; // sw $fp $t5 6
		  memoria_hd[368] = 32'b00001111101001100000000000000101; // lw $fp $t6 5
		  memoria_hd[369] = 32'b00000100110001100000000000000000; // addi $t6 $t6 0
		  memoria_hd[370] = 32'b00010011101001100000000000000101; // sw $fp $t6 5
		  memoria_hd[371] = 32'b00000100000110110000000000000000; // addi $aux $zero 0
		  memoria_hd[372] = 32'b00000000101110110011100000000001; // sub $t7 $t5 $aux
		  memoria_hd[373] = 32'b00011000000001110000000000011011; // bne $t7 $zero 27
		  memoria_hd[374] = 32'b00001111101010000000000000000011; // lw $fp $t8 3
		  memoria_hd[375] = 32'b00000101000111000000000000000000; // addi $gp $t8 0
		  memoria_hd[376] = 32'b00011100000000000000000000110100; // jump 52
		  memoria_hd[377] = 32'b00000000101000010100100000100100; // sle $t9 $t5 $t1
		  memoria_hd[378] = 32'b00010100000010010000000000110011; // beq $t9 $zero 51
		  memoria_hd[379] = 32'b00001111101010100000000000000101; // lw $fp $t10 5
		  memoria_hd[380] = 32'b00001111101010110000000000000011; // lw $fp $t11 3
		  memoria_hd[381] = 32'b00001111101011000000000000000100; // lw $fp $t12 4
		  memoria_hd[382] = 32'b00000001011011000110100000000000; // add $t13 $t11 $t12
		  memoria_hd[383] = 32'b00000101101010100000000000000000; // addi $t10 $t13 0
		  memoria_hd[384] = 32'b00010011101010100000000000000101; // sw $fp $t10 5
		  memoria_hd[385] = 32'b00001111101011100000000000000011; // lw $fp $t14 3
		  memoria_hd[386] = 32'b00001111101011110000000000000100; // lw $fp $t15 4
		  memoria_hd[387] = 32'b00000101111011100000000000000000; // addi $t14 $t15 0
		  memoria_hd[388] = 32'b00010011101011100000000000000011; // sw $fp $t14 3
		  memoria_hd[389] = 32'b00001111101100000000000000000100; // lw $fp $t16 4
		  memoria_hd[390] = 32'b00001111101100010000000000000101; // lw $fp $t17 5
		  memoria_hd[391] = 32'b00000110001100000000000000000000; // addi $t16 $t17 0
		  memoria_hd[392] = 32'b00010011101100000000000000000100; // sw $fp $t16 4
		  memoria_hd[393] = 32'b00001111101100100000000000000110; // lw $fp $t18 6
		  memoria_hd[394] = 32'b00001111101100110000000000000110; // lw $fp $t19 6
		  memoria_hd[395] = 32'b00000100000110110000000000000001; // addi $aux $zero 1
		  memoria_hd[396] = 32'b00000010011110111010000000000000; // add $t20 $t19 $aux
		  memoria_hd[397] = 32'b00000110100100100000000000000000; // addi $t18 $t20 0
		  memoria_hd[398] = 32'b00010011101100100000000000000110; // sw $fp $t18 6
		  memoria_hd[399] = 32'b00000110100001010000000000000000; // addi $t5 $t20 0
		  memoria_hd[400] = 32'b00011100000000000000000000011011; // jump 27
		  memoria_hd[401] = 32'b00011100000000000000000000110100; // jump 52
		  memoria_hd[402] = 32'b00001111101101010000000000000100; // lw $fp $t21 4
		  memoria_hd[403] = 32'b00000110101111000000000000000000; // addi $gp $t21 0
		  memoria_hd[404] = 32'b00001111101111110000000000000001; // lw $fp $ra 1
		  memoria_hd[405] = 32'b00100111111000000000000000000000; // jr $ra $zero $zero
		  memoria_hd[406] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[407] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[408] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[409] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[410] = 32'b00101100000000101111111111111111; // input $t2
		  memoria_hd[411] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[412] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[413] = 32'b00001111101000110000000000000000; // lw $fp $t3 0
		  memoria_hd[414] = 32'b00010011110111010000000000000000; // sw $sp $fp 0
		  memoria_hd[415] = 32'b00000111110111010000000000000000; // addi $fp $sp 0
		  memoria_hd[416] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[417] = 32'b00010011101000110000000000000010; // sw $fp $t3 2
		  memoria_hd[418] = 32'b00110000000000000000000000000001; // jal 1
		  memoria_hd[419] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[420] = 32'b00001111101111010000000000000000; // lw $fp $fp 0
		  memoria_hd[421] = 32'b00000111100001000000000000000000; // addi $t4 $gp 0
		  memoria_hd[422] = 32'b00101000100111111111111111111111; // output $t4
		  memoria_hd[423] = 32'b11111000000000000000000000000000; // halt 
		  
		  // Programa 3 - Calcula 
		  /*memoria_hd[500] = 32'b00011100000000000000000000010010; // jump 18 
		  memoria_hd[501] = 32'b00010011101111110000000000000001; // sw $fp $ra 1
		  memoria_hd[502] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[503] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[504] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[505] = 32'b00001111101000010000000000000010; // lw $fp $t1 2
		  memoria_hd[506] = 32'b00001111101000100000000000000011; // lw $fp $t2 3
		  memoria_hd[507] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[508] = 32'b00001111101001000000000000000100; // lw $fp $t4 4
		  memoria_hd[509] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[510] = 32'b00001111101001100000000000000011; // lw $fp $t6 3
		  memoria_hd[511] = 32'b00000000101001100011100000000000; // add $t7 $t5 $t6
		  memoria_hd[512] = 32'b00000100111001000000000000000000; // addi $t4 $t7 0
		  memoria_hd[513] = 32'b00010011101001000000000000000100; // sw $fp $t4 4
		  memoria_hd[514] = 32'b00001111101010000000000000000100; // lw $fp $t8 4
		  memoria_hd[515] = 32'b00000101000111000000000000000000; // addi $gp $t8 0
		  memoria_hd[516] = 32'b00001111101111110000000000000001; // lw $fp $ra 1
		  memoria_hd[517] = 32'b00100111111000000000000000000000; // jr $ra $zero $zero
		  memoria_hd[518] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[519] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[520] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[521] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[522] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[523] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[524] = 32'b00101100000000101111111111111111; // input $t2
		  memoria_hd[525] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0  
		  memoria_hd[526] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[527] = 32'b00001111101000110000000000000001; // lw $fp $t3 1
		  memoria_hd[528] = 32'b00101100000001001111111111111111; // input $t4  
		  memoria_hd[529] = 32'b00000100100000110000000000000000; // addi $t3 $t4 0
		  memoria_hd[530] = 32'b00010011101000110000000000000001; // sw $fp $t3 1
		  memoria_hd[531] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[532] = 32'b00001111101001100000000000000000; // lw $fp $t6 0
		  memoria_hd[533] = 32'b00001111101001110000000000000001; // lw $fp $t7 1
		  memoria_hd[534] = 32'b00010011110111010000000000000000; // sw $sp $fp 0
		  memoria_hd[535] = 32'b00000111110111010000000000000000; // addi $fp $sp 0
		  memoria_hd[536] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[537] = 32'b00010011101001110000000000000011; // sw $fp $t7 3
		  memoria_hd[538] = 32'b00010011101001100000000000000010; // sw $fp $t6 2
		  memoria_hd[539] = 32'b00110000000000000000000000000001; // jal 1
		  memoria_hd[540] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[541] = 32'b00001111101111010000000000000000; // lw $fp $fp 0
		  memoria_hd[542] = 32'b00000111100010000000000000000000; // addi $t8 $gp 0
		  memoria_hd[543] = 32'b00000101000001010000000000000000; // addi $t5 $t8 0
		  memoria_hd[544] = 32'b00010011101001010000000000000010; // sw $fp $t5 2
		  memoria_hd[545] = 32'b00001111101010010000000000000010; // lw $fp $t9 2
		  memoria_hd[546] = 32'b00101001001111111111111111111111; // output $t9  
		  memoria_hd[547] = 32'b11111000000000000000000000000000; // halt*/

		  memoria_hd[500] = 32'b00011100000000000000000000000001; // jump 1 
		  memoria_hd[501] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[502] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[503] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[504] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[505] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[506] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[507] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[508] = 32'b00101100000000101111111111111111; // input $t2
		  memoria_hd[509] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[510] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[511] = 32'b00001111101000110000000000000001; // lw $fp $t3 1
		  memoria_hd[512] = 32'b00101100000001001111111111111111; // input $t4
		  memoria_hd[513] = 32'b00000100100000110000000000000000; // addi $t3 $t4 0
		  memoria_hd[514] = 32'b00010011101000110000000000000001; // sw $fp $t3 1
		  memoria_hd[515] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[516] = 32'b00001111101001100000000000000000; // lw $fp $t6 0
		  memoria_hd[517] = 32'b00001111101001110000000000000001; // lw $fp $t7 1
		  memoria_hd[518] = 32'b00000000110001110100000000000010; // mult $t8 $t6 $t7
		  memoria_hd[519] = 32'b00000101000001010000000000000000; // addi $t5 $t8 0
		  memoria_hd[520] = 32'b00010011101001010000000000000010; // sw $fp $t5 2
		  memoria_hd[521] = 32'b00001111101010010000000000000011; // lw $fp $t9 3
		  memoria_hd[522] = 32'b00101100000010101111111111111111; // input $t10 
		  memoria_hd[523] = 32'b00000101010010010000000000000000; // addi $t9 $t10 0
		  memoria_hd[524] = 32'b00010011101010010000000000000011; // sw $fp $t9 3
		  memoria_hd[525] = 32'b00001111101010110000000000000010; // lw $fp $t11 2
		  memoria_hd[526] = 32'b00001111101011000000000000000010; // lw $fp $t12 2
		  memoria_hd[527] = 32'b00001111101011010000000000000011; // lw $fp $t13 3
		  memoria_hd[528] = 32'b00000001100011010111000000000001; // sub $t14 $t12 $t13
		  memoria_hd[529] = 32'b00000101110010110000000000000000; // addi $t11 $t14 0
		  memoria_hd[530] = 32'b00010011101010110000000000000010; // sw $fp $t11 2
		  memoria_hd[531] = 32'b00001111101011110000000000000010; // lw $fp $t15 2
		  memoria_hd[532] = 32'b00101001111111111111111111111111; // output $t15
		  memoria_hd[533] = 32'b11111000000000000000000000000000; // halt


		  
		  // Programa 4 - Potencia 
		  memoria_hd[650] = 32'b00011100000000000000000000100011; // jump 35 
		  memoria_hd[651] = 32'b00010011101111110000000000000001; // sw $fp $ra 1
		  memoria_hd[652] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[653] = 32'b00000111110111100000000000000001; // addi $sp $sp 1 
		  memoria_hd[654] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[655] = 32'b00001111101000010000000000000010; // lw $fp $t1 2
		  memoria_hd[656] = 32'b00001111101000100000000000000011; // lw $fp $t2 3
		  memoria_hd[657] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[658] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[659] = 32'b00001111101001000000000000000101; // lw $fp $t4 5
		  memoria_hd[660] = 32'b00000100100001000000000000000001; // addi $t4 $t4 1
		  memoria_hd[661] = 32'b00010011101001000000000000000101; // sw $fp $t4 5
		  memoria_hd[662] = 32'b00001111101001010000000000000100; // lw $fp $t5 4
		  memoria_hd[663] = 32'b00000100101001010000000000000000; // addi $t5 $t5 0
		  memoria_hd[664] = 32'b00010011101001010000000000000100; // sw $fp $t5 4
		  memoria_hd[665] = 32'b00000000101000100011000000000111; // slt $t6 $t5 $t2
		  memoria_hd[666] = 32'b00010100000001100000000000011111; // beq $t6 $zero 31
		  memoria_hd[667] = 32'b00001111101001110000000000000101; // lw $fp $t7 5
		  memoria_hd[668] = 32'b00001111101010000000000000000101; // lw $fp $t8 5
		  memoria_hd[669] = 32'b00001111101010010000000000000010; // lw $fp $t9 2
		  memoria_hd[670] = 32'b00000001000010010101000000000010; // mult $t10 $t8 $t9
		  memoria_hd[671] = 32'b00000101010001110000000000000000; // addi $t7 $t10 0
		  memoria_hd[672] = 32'b00010011101001110000000000000101; // sw $fp $t7 5
		  memoria_hd[673] = 32'b00001111101010110000000000000011; // lw $fp $t11 3
		  memoria_hd[674] = 32'b00001111101011000000000000000011; // lw $fp $t12 3
		  memoria_hd[675] = 32'b00000100000110110000000000000001; // addi $aux $zero 1
		  memoria_hd[676] = 32'b00000001100110110110100000000001; // sub $t13 $t12 $aux
		  memoria_hd[677] = 32'b00000101101010110000000000000000; // addi $t11 $t13 0
		  memoria_hd[678] = 32'b00010011101010110000000000000011; // sw $fp $t11 3
		  memoria_hd[679] = 32'b00000101101000100000000000000000; // addi $t2 $t13 0
		  memoria_hd[680] = 32'b00011100000000000000000000001111; // jump 15
		  memoria_hd[681] = 32'b00001111101011100000000000000101; // lw $fp $t14 5
		  memoria_hd[682] = 32'b00000101110111000000000000000000; // addi $gp $t14 0
		  memoria_hd[683] = 32'b00001111101111110000000000000001; // lw $fp $ra 1
		  memoria_hd[684] = 32'b00100111111000000000000000000000; // jr $ra $zero $zero
		  memoria_hd[685] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[686] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[687] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[688] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[689] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[690] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[691] = 32'b00101100000000101111111111111111; // input $t2
		  memoria_hd[692] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[693] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[694] = 32'b00001111101000110000000000000001; // lw $fp $t3 1
		  memoria_hd[695] = 32'b00101100000001001111111111111111; // input $t4 
		  memoria_hd[696] = 32'b00000100100000110000000000000000; // addi $t3 $t4 0
		  memoria_hd[697] = 32'b00010011101000110000000000000001; // sw $fp $t3 1
		  memoria_hd[698] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[699] = 32'b00001111101001100000000000000000; // lw $fp $t6 0
		  memoria_hd[700] = 32'b00001111101001110000000000000001; // lw $fp $t7 1
		  memoria_hd[701] = 32'b00010011110111010000000000000000; // sw $sp $fp 0
		  memoria_hd[702] = 32'b00000111110111010000000000000000; // addi $fp $sp 0
		  memoria_hd[703] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[704] = 32'b00010011101001110000000000000011; // sw $fp $t7 3
		  memoria_hd[705] = 32'b00010011101001100000000000000010; // sw $fp $t6 2
		  memoria_hd[706] = 32'b00110000000000000000000000000001; // jal 1
		  memoria_hd[707] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[708] = 32'b00001111101111010000000000000000; // lw $fp $fp 0
		  memoria_hd[709] = 32'b00000111100010000000000000000000; // addi $t8 $gp 0
		  memoria_hd[710] = 32'b00000101000001010000000000000000; // addi $t5 $t8 0
		  memoria_hd[711] = 32'b00010011101001010000000000000010; // sw $fp $t5 2
		  memoria_hd[712] = 32'b00001111101010010000000000000010; // lw $fp $t9 2
		  memoria_hd[713] = 32'b00101001001111111111111111111111; // output $t9
		  memoria_hd[714] = 32'b11111000000000000000000000000000; // halt
		  
		  // Programa 5 - Media 
		  memoria_hd[800] = 32'b00011100000000000000000000000001; // jump 1  
		  memoria_hd[801] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[802] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[803] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[804] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[805] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[806] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[807] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[808] = 32'b00101100000000101111111111111111; // input $t2
		  memoria_hd[809] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[810] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[811] = 32'b00001111101000110000000000000001; // lw $fp $t3 1
		  memoria_hd[812] = 32'b00101100000001001111111111111111; // input $t4
		  memoria_hd[813] = 32'b00000100100000110000000000000000; // addi $t3 $t4 0
		  memoria_hd[814] = 32'b00010011101000110000000000000001; // sw $fp $t3 1
		  memoria_hd[815] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[816] = 32'b00101100000001101111111111111111; // input $t6
		  memoria_hd[817] = 32'b00000100110001010000000000000000; // addi $t5 $t6 0
		  memoria_hd[818] = 32'b00010011101001010000000000000010; // sw $fp $t5 2
		  memoria_hd[819] = 32'b00001111101001110000000000000011; // lw $fp $t7 3
		  memoria_hd[820] = 32'b00001111101010000000000000000000; // lw $fp $t8 0
		  memoria_hd[821] = 32'b00001111101010010000000000000001; // lw $fp $t9 1
		  memoria_hd[822] = 32'b00000001000010010101000000000000; // add $t10 $t8 $t9
		  memoria_hd[823] = 32'b00001111101010110000000000000010; // lw $fp $t11 2
		  memoria_hd[824] = 32'b00000001010010110110000000000000; // add $t12 $t10 $t11
		  memoria_hd[825] = 32'b00000100000110110000000000000011; // addi $aux $zero 3
		  memoria_hd[826] = 32'b00000001100110110110100000000011; // div $t13 $t12 $aux
		  memoria_hd[827] = 32'b00000101101001110000000000000000; // addi $t7 $t13 0
		  memoria_hd[828] = 32'b00010011101001110000000000000011; // sw $fp $t7 3
		  memoria_hd[829] = 32'b00001111101011100000000000000011; // lw $fp $t14 3
		  memoria_hd[830] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[831] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[832] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[833] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[835] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[836] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[837] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[838] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[839] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[840] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[841] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[842] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[843] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[844] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[845] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[846] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[847] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[848] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[849] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[850] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[851] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[852] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[853] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[854] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[855] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[856] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[857] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[858] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[859] = 32'b00110100000000000000000000000000; // nop
		  memoria_hd[860] = 32'b00101001110111111111111111111111; // output $t14
		  memoria_hd[861] = 32'b11111000000000000000000000000000; // halt
		  
		  // Programa 6 - Área triângulo 
		  memoria_hd[950] = 32'b00011100000000000000000000000001; // jump 1
		  memoria_hd[951] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[952] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[953] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[954] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[955] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[956] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[957] = 32'b00101100000000101111111111111111; // input $t2
		  memoria_hd[958] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[959] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[960] = 32'b00001111101000110000000000000001; // lw $fp $t3 1
		  memoria_hd[961] = 32'b00101100000001001111111111111111; // input $t4
		  memoria_hd[962] = 32'b00000100100000110000000000000000; // addi $t3 $t4 0
		  memoria_hd[963] = 32'b00010011101000110000000000000001; // sw $fp $t3 1
		  memoria_hd[964] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[965] = 32'b00001111101001100000000000000000; // lw $fp $t6 0
		  memoria_hd[966] = 32'b00001111101001110000000000000001; // lw $fp $t7 1
		  memoria_hd[967] = 32'b00000000110001110100000000000010; // mult $t8 $t6 $t7
		  memoria_hd[968] = 32'b00000100000110110000000000000010; // addi $aux $zero 2
		  memoria_hd[969] = 32'b00000001000110110100100000000011; // div $t9 $t8 $aux
		  memoria_hd[970] = 32'b00000101001001010000000000000000; // addi $t5 $t9 0
		  memoria_hd[971] = 32'b00010011101001010000000000000010; // sw $fp $t5 2
		  memoria_hd[972] = 32'b00001111101010100000000000000010; // lw $fp $t10 2
		  memoria_hd[973] = 32'b00101001010111111111111111111111; // output $t10
		  memoria_hd[974] = 32'b11111000000000000000000000000000; // halt
		  
		  // Programa 7 - Fatorial 
		  memoria_hd[1100] = 32'b00011100000000000000000000100111; // jump 39	  
		  memoria_hd[1101] = 32'b00010011101111110000000000000001; // sw $fp $ra 1
		  memoria_hd[1102] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1103] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1104] = 32'b00001111101000010000000000000010; // lw $fp $t1 2
		  memoria_hd[1105] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1106] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1107] = 32'b00000100000110110000000000000001; // addi $aux $zero 1
		  memoria_hd[1108] = 32'b00000000001110110001100000000001; // sub $t3 $t1 $aux
		  memoria_hd[1109] = 32'b00011000000000110000000000001100; // bne $t3 $zero 12
		  memoria_hd[1110] = 32'b00000111100111000000000000000001; // addi $gp $gp 1
		  memoria_hd[1111] = 32'b00011100000000000000000000100101; // jump 37
		  memoria_hd[1112] = 32'b00001111101001000000000000000100; // lw $fp $t4 4
		  memoria_hd[1113] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[1114] = 32'b00000100000110110000000000000001; // addi $aux $zero 1
		  memoria_hd[1115] = 32'b00000000101110110011000000000001; // sub $t6 $t5 $aux
		  memoria_hd[1116] = 32'b00000100110001000000000000000000; // addi $t4 $t6 0
		  memoria_hd[1117] = 32'b00010011101001000000000000000100; // sw $fp $t4 4
		  memoria_hd[1118] = 32'b00001111101001110000000000000011; // lw $fp $t7 3
		  memoria_hd[1119] = 32'b00001111101010000000000000000010; // lw $fp $t8 2
		  memoria_hd[1120] = 32'b00010011101010000000000000110010; // sw $fp $t8 50
		  memoria_hd[1121] = 32'b00001111101010010000000000000100; // lw $fp $t9 4
		  memoria_hd[1122] = 32'b00010011110111010000000000000000; // sw $sp $fp 0
		  memoria_hd[1123] = 32'b00000111110111010000000000000000; // addi $fp $sp 0
		  memoria_hd[1124] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1125] = 32'b00010011101010010000000000000010; // sw $fp $t9 2
		  memoria_hd[1126] = 32'b00110000000000000000000000000001; // jal 1
		  memoria_hd[1127] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[1128] = 32'b00001111101111010000000000000000; // lw $fp $fp 0
		  memoria_hd[1129] = 32'b00000111100010100000000000000000; // addi $t10 $gp 0
		  memoria_hd[1130] = 32'b00001111101010000000000000110010; // lw $fp $t8 50
		  memoria_hd[1131] = 32'b00000001000010100101100000000010; // mult $t11 $t8 $t10
		  memoria_hd[1132] = 32'b00000101011001110000000000000000; // addi $t7 $t11 0
		  memoria_hd[1133] = 32'b00010011101001110000000000000011; // sw $fp $t7 3
		  memoria_hd[1134] = 32'b00001111101011000000000000000011; // lw $fp $t12 3
		  memoria_hd[1135] = 32'b00000101100111000000000000000000; // addi $gp $t12 0
		  memoria_hd[1136] = 32'b00011100000000000000000000100101; // jump 37
		  memoria_hd[1137] = 32'b00001111101111110000000000000001; // lw $fp $ra 1
		  memoria_hd[1138] = 32'b00100111111000000000000000000000; // jr $ra $zero $zero
		  memoria_hd[1139] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[1140] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[1141] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1142] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1143] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[1144] = 32'b00101100000000101111111111111111; // input $t2  
		  memoria_hd[1145] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[1146] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[1147] = 32'b00001111101000110000000000000001; // lw $fp $t3 1
		  memoria_hd[1148] = 32'b00001111101001000000000000000000; // lw $fp $t4 0
		  memoria_hd[1149] = 32'b00010011110111010000000000000000; // sw $sp $fp 0
		  memoria_hd[1150] = 32'b00000111110111010000000000000000; // addi $fp $sp 0
		  memoria_hd[1151] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1152] = 32'b00010011101001000000000000000010; // sw $fp $t4 2
		  memoria_hd[1153] = 32'b00110000000000000000000000000001; // jal 1
		  memoria_hd[1154] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[1155] = 32'b00001111101111010000000000000000; // lw $fp $fp 0
		  memoria_hd[1156] = 32'b00000111100001010000000000000000; // addi $t5 $gp 0
		  memoria_hd[1157] = 32'b00000100101000110000000000000000; // addi $t3 $t5 0
		  memoria_hd[1158] = 32'b00010011101000110000000000000001; // sw $fp $t3 1
		  memoria_hd[1159] = 32'b00001111101001100000000000000001; // lw $fp $t6 1
		  memoria_hd[1160] = 32'b00101000110111111111111111111111; // output $t6 
		  memoria_hd[1161] = 32'b11111000000000000000000000000000; // halt
		  
		  // Programa 8 - Contagem regressiva 
		  memoria_hd[1250] = 32'b00011100000000000000000000000001; // jump 1
		  memoria_hd[1251] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[1252] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[1253] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1254] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1255] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[1256] = 32'b00101100000000101111111111111111; // input $t2 
		  memoria_hd[1257] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[1258] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[1259] = 32'b00000100000110110000000000000000; // addi $aux $zero 0
		  memoria_hd[1260] = 32'b00000011011000010001100000000111; // slt $t3 $aux $t1
		  memoria_hd[1261] = 32'b00010100000000110000000000011010; // beq $t3 $zero 26
		  memoria_hd[1262] = 32'b00001111101001000000000000000000; // lw $fp $t4 0
		  memoria_hd[1263] = 32'b00101000100111111111111111111111; // output $t4
		  memoria_hd[1264] = 32'b00001111101001100000000000000001; // lw $fp $t6 1
		  memoria_hd[1265] = 32'b00101100000001111111111111111111; // input $t7  
		  memoria_hd[1266] = 32'b00000100111001100000000000000000; // addi $t6 $t7 0
		  memoria_hd[1267] = 32'b00010011101001100000000000000001; // sw $fp $t6 1
		  memoria_hd[1268] = 32'b00001111101010000000000000000000; // lw $fp $t8 0
		  memoria_hd[1269] = 32'b00001111101010010000000000000000; // lw $fp $t9 0
		  memoria_hd[1270] = 32'b00000100000110110000000000000001; // addi $aux $zero 1
		  memoria_hd[1271] = 32'b00000001001110110101000000000001; // sub $t10 $t9 $aux
		  memoria_hd[1272] = 32'b00000101010010000000000000000000; // addi $t8 $t10 0
		  memoria_hd[1273] = 32'b00010011101010000000000000000000; // sw $fp $t8 0
		  memoria_hd[1274] = 32'b00000101010000010000000000000000; // addi $t1 $t10 0
		  memoria_hd[1275] = 32'b00011100000000000000000000001001; // jump 9 
		  memoria_hd[1276] = 32'b11111000000000000000000000000000; // halt
		  
		  // Programa 9 - Calculadora  
		  memoria_hd[1400] = 32'b00011100000000000000000000000001; // jump 1
		  memoria_hd[1401] = 32'b00000100000111010000000000111100; // addi $fp $zero 60
		  memoria_hd[1402] = 32'b00000111101111100000000000000000; // addi $sp $fp 0
		  memoria_hd[1403] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1404] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1405] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1406] = 32'b00000111110111100000000000000001; // addi $sp $sp 1
		  memoria_hd[1407] = 32'b00001111101000010000000000000000; // lw $fp $t1 0
		  memoria_hd[1408] = 32'b00101100000000101111111111111111; // input $t2 
		  memoria_hd[1409] = 32'b00000100010000010000000000000000; // addi $t1 $t2 0
		  memoria_hd[1410] = 32'b00010011101000010000000000000000; // sw $fp $t1 0
		  memoria_hd[1411] = 32'b00001111101000110000000000000001; // lw $fp $t3 1
		  memoria_hd[1412] = 32'b00101100000001001111111111111111; // input $t4
		  memoria_hd[1413] = 32'b00000100100000110000000000000000; // addi $t3 $t4 0
		  memoria_hd[1414] = 32'b00010011101000110000000000000001; // sw $fp $t3 1
		  memoria_hd[1415] = 32'b00001111101001010000000000000010; // lw $fp $t5 2
		  memoria_hd[1416] = 32'b00101100000001101111111111111111; // input $t6
		  memoria_hd[1417] = 32'b00000100110001010000000000000000; // addi $t5 $t6 0
		  memoria_hd[1418] = 32'b00010011101001010000000000000010; // sw $fp $t5 2
		  memoria_hd[1419] = 32'b00000100000110110000000000000001; // addi $aux $zero 1
		  memoria_hd[1420] = 32'b00000000001110110011100000000001; // sub $t7 $t1 $aux
		  memoria_hd[1421] = 32'b00011000000001110000000000011101; // bne $t7 $zero 29
		  memoria_hd[1422] = 32'b00001111101010000000000000000011; // lw $fp $t8 3
		  memoria_hd[1423] = 32'b00001111101010010000000000000001; // lw $fp $t9 1
		  memoria_hd[1424] = 32'b00001111101010100000000000000010; // lw $fp $t10 2
		  memoria_hd[1425] = 32'b00000001001010100101100000000000; // add $t11 $t9 $t10
		  memoria_hd[1426] = 32'b00000101011010000000000000000000; // addi $t8 $t11 0
		  memoria_hd[1427] = 32'b00010011101010000000000000000011; // sw $fp $t8 3
		  memoria_hd[1428] = 32'b00011100000000000000000000111010; // jump 58
		  memoria_hd[1429] = 32'b00000100000110110000000000000010; // addi $aux $zero 2
		  memoria_hd[1430] = 32'b00000000001110110110000000000001; // sub $t12 $t1 $aux
		  memoria_hd[1431] = 32'b00011000000011000000000000100111; // bne $t12 $zero 39
		  memoria_hd[1432] = 32'b00001111101011010000000000000011; // lw $fp $t13 3
		  memoria_hd[1433] = 32'b00001111101011100000000000000001; // lw $fp $t14 1
		  memoria_hd[1434] = 32'b00001111101011110000000000000010; // lw $fp $t15 2
		  memoria_hd[1435] = 32'b00000001110011111000000000000001; // sub $t16 $t14 $t15
		  memoria_hd[1436] = 32'b00000110000011010000000000000000; // addi $t13 $t16 0
		  memoria_hd[1437] = 32'b00010011101011010000000000000011; // sw $fp $t13 3
		  memoria_hd[1438] = 32'b00011100000000000000000000111001; // jump 57 
		  memoria_hd[1439] = 32'b00000100000110110000000000000011; // addi $aux $zero 3
		  memoria_hd[1440] = 32'b00000000001110111000100000000001; // sub $t17 $t1 $aux
		  memoria_hd[1441] = 32'b00011000000100010000000000110001; // bne $t17 $zero 49
		  memoria_hd[1442] = 32'b00001111101100100000000000000011; // lw $fp $t18 3
		  memoria_hd[1443] = 32'b00001111101100110000000000000001; // lw $fp $t19 1
		  memoria_hd[1444] = 32'b00001111101101000000000000000010; // lw $fp $t20 2
		  memoria_hd[1445] = 32'b00000010011101001010100000000010; // mult $t21 $t19 $t20
	     memoria_hd[1446] = 32'b00000110101100100000000000000000; // addi $t18 $t21 0
	     memoria_hd[1447] = 32'b00010011101100100000000000000011; // sw $fp $t18 3
		  memoria_hd[1448] = 32'b00011100000000000000000000111000; // jump 56
		  memoria_hd[1449] = 32'b00001111101101100000000000000011; // lw $fp $t22 3
		  memoria_hd[1450] = 32'b00001111101101110000000000000001; // lw $fp $t23 1
		  memoria_hd[1451] = 32'b00001111101110000000000000000010; // lw $fp $t24 2
		  memoria_hd[1452] = 32'b00000010111110001100100000000011; // div $t25 $t23 $t24
		  memoria_hd[1453] = 32'b00000111001101100000000000000000; // addi $t22 $t25 0
		  memoria_hd[1454] = 32'b00010011101101100000000000000011; // sw $fp $t22 3
		  memoria_hd[1455] = 32'b00011100000000000000000000111000; // jump 56
		  memoria_hd[1456] = 32'b00011100000000000000000000111001; // jump 57
		  memoria_hd[1457] = 32'b00011100000000000000000000111010; // jump 58
		  memoria_hd[1458] = 32'b00001111101110100000000000000011; // lw $fp $t26 3
		  memoria_hd[1459] = 32'b00101011010111111111111111111111; // output $t26
		  memoria_hd[1460] = 32'b11111000000000000000000000000000; // halt
		  
		  /*// Programa 10 - Maior  
		  memoria_hd[1550] = 32'b00011100000000000000000000000001; // jump 1*/
		  
		  
    end

    always @(posedge Clock) begin
        instrucao <= memoria_hd[addr];
    end
endmodule